`define READ_VALID 1'b1
`define WRITE_VALID 1'b0

`define FULL 1'b1
`define EMPTY 1'b0

module ProgramCache (clk, addr, data_out);
    input clk;
	input [9:0] addr;

    output [31:0] data_out;
	//2**32-1 = 4,294,967,295
    reg [7:0] data[1023:0];

	assign data_out = {data[addr], data[addr+1], data[addr+2], data[addr+3]};

    initial begin
		// 188225285 ADD -575174121 = -386948836
		//H 0b381705 ADD a24875e9 = 97105ee4
		data[0] = 8'b00111100;
		data[1] = 8'b00000001;
		data[2] = 8'b00001011;
		data[3] = 8'b00111000;
		data[4] = 8'b00110100;
		data[5] = 8'b00100001;
		data[6] = 8'b00010111;
		data[7] = 8'b00000101;
		data[8] = 8'b00111100;
		data[9] = 8'b00000010;
		data[10] = 8'b10100010;
		data[11] = 8'b01001000;
		data[12] = 8'b00110100;
		data[13] = 8'b01000010;
		data[14] = 8'b01110101;
		data[15] = 8'b11101001;
		data[16] = 8'b00000000;
		data[17] = 8'b00100010;
		data[18] = 8'b11111000;
		data[19] = 8'b00100000;
		// -606441343 ADDI 26006 = -606415337
		//H a4258f7f ADDI 00006596 = a42529e9
		data[20] = 8'b00111100;
		data[21] = 8'b00000001;
		data[22] = 8'b10100100;
		data[23] = 8'b00100101;
		data[24] = 8'b00110100;
		data[25] = 8'b00100001;
		data[26] = 8'b10001111;
		data[27] = 8'b01111111;
		data[28] = 8'b00100000;
		data[29] = 8'b00111111;
		data[30] = 8'b01100101;
		data[31] = 8'b10010110;
		// 4254819324 ADDU 1558667430 = 5813486754
		//H fd9b63fc ADDU 5ce760a6 = 0x1_5a82c4a2
		data[32] = 8'b00111100;
		data[33] = 8'b00000001;
		data[34] = 8'b11111101;
		data[35] = 8'b10011011;
		data[36] = 8'b00110100;
		data[37] = 8'b00100001;
		data[38] = 8'b01100011;
		data[39] = 8'b11111100;
		data[40] = 8'b00111100;
		data[41] = 8'b00000010;
		data[42] = 8'b01011100;
		data[43] = 8'b11100111;
		data[44] = 8'b00110100;
		data[45] = 8'b01000010;
		data[46] = 8'b01100000;
		data[47] = 8'b10100110;
		data[48] = 8'b00000000;
		data[49] = 8'b00100010;
		data[50] = 8'b11111000;
		data[51] = 8'b00100001;
		// -1680872635 ADDIU 24663 = -1680847972
		//H e43014bb ADDIU 00006057 = e42fb464
		data[52] = 8'b00111100;
		data[53] = 8'b00000001;
		data[54] = 8'b11100100;
		data[55] = 8'b00110000;
		data[56] = 8'b00110100;
		data[57] = 8'b00100001;
		data[58] = 8'b00010100;
		data[59] = 8'b10111011;
		data[60] = 8'b00100100;
		data[61] = 8'b00111111;
		data[62] = 8'b01100000;
		data[63] = 8'b01010111;
		// 547813419 SUB 228591612 = 319221807
		//H 20a6f82b SUB 0da007fc = 1306f02f
		data[64] = 8'b00111100;
		data[65] = 8'b00000001;
		data[66] = 8'b00100000;
		data[67] = 8'b10100110;
		data[68] = 8'b00110100;
		data[69] = 8'b00100001;
		data[70] = 8'b11111000;
		data[71] = 8'b00101011;
		data[72] = 8'b00111100;
		data[73] = 8'b00000010;
		data[74] = 8'b00001101;
		data[75] = 8'b10100000;
		data[76] = 8'b00110100;
		data[77] = 8'b01000010;
		data[78] = 8'b00000111;
		data[79] = 8'b11111100;
		data[80] = 8'b00000000;
		data[81] = 8'b00100010;
		data[82] = 8'b11111000;
		data[83] = 8'b00100010;
		// 2063490976 SLT -1546272794 = False
		//H 7afe5fa0 SLT dc2a401a = 00000000
		data[84] = 8'b00111100;
		data[85] = 8'b00000001;
		data[86] = 8'b01111010;
		data[87] = 8'b11111110;
		data[88] = 8'b00110100;
		data[89] = 8'b00100001;
		data[90] = 8'b01011111;
		data[91] = 8'b10100000;
		data[92] = 8'b00111100;
		data[93] = 8'b00000010;
		data[94] = 8'b11011100;
		data[95] = 8'b00101010;
		data[96] = 8'b00110100;
		data[97] = 8'b01000010;
		data[98] = 8'b01000000;
		data[99] = 8'b00011010;
		data[100] = 8'b00000000;
		data[101] = 8'b00100010;
		data[102] = 8'b11111000;
		data[103] = 8'b00101010;
		// -2026551683 MUL 1915526345 = -3881913138290588635
		//H f8cab983 MUL 722c9cc9 = 67448424
		data[104] = 8'b00111100;
		data[105] = 8'b00000001;
		data[106] = 8'b11111000;
		data[107] = 8'b11001010;
		data[108] = 8'b00110100;
		data[109] = 8'b00100001;
		data[110] = 8'b10111001;
		data[111] = 8'b10000011;
		data[112] = 8'b00111100;
		data[113] = 8'b00000010;
		data[114] = 8'b01110010;
		data[115] = 8'b00101100;
		data[116] = 8'b00110100;
		data[117] = 8'b01000010;
		data[118] = 8'b10011100;
		data[119] = 8'b11001001;
		data[120] = 8'b01110000;
		data[121] = 8'b00100010;
		data[122] = 8'b11111000;
		data[123] = 8'b00000010;
		// 3378638932 AND 1682394321 = 1078018128
		//H c961f054 AND 64474cd1 = 40414050
		data[124] = 8'b00111100;
		data[125] = 8'b00000001;
		data[126] = 8'b11001001;
		data[127] = 8'b01100001;
		data[128] = 8'b00110100;
		data[129] = 8'b00100001;
		data[130] = 8'b11110000;
		data[131] = 8'b01010100;
		data[132] = 8'b00111100;
		data[133] = 8'b00000010;
		data[134] = 8'b01100100;
		data[135] = 8'b01000111;
		data[136] = 8'b00110100;
		data[137] = 8'b01000010;
		data[138] = 8'b01001100;
		data[139] = 8'b11010001;
		data[140] = 8'b00000000;
		data[141] = 8'b00100010;
		data[142] = 8'b11111000;
		data[143] = 8'b00100100;
		// 1800125538 ANDI 45566 = 45154
		//H 6b4bbc62 ANDI 0000b1fe = 0000b062
		data[144] = 8'b00111100;
		data[145] = 8'b00000001;
		data[146] = 8'b01101011;
		data[147] = 8'b01001011;
		data[148] = 8'b00110100;
		data[149] = 8'b00100001;
		data[150] = 8'b10111100;
		data[151] = 8'b01100010;
		data[152] = 8'b00110000;
		data[153] = 8'b00111111;
		data[154] = 8'b10110001;
		data[155] = 8'b11111110;
		// 1679827541 OR 1590071485 = 2129048317
		//H 64202255 OR 5ec690bd = 7ee6b2fd
		data[156] = 8'b00111100;
		data[157] = 8'b00000001;
		data[158] = 8'b01100100;
		data[159] = 8'b00100000;
		data[160] = 8'b00110100;
		data[161] = 8'b00100001;
		data[162] = 8'b00100010;
		data[163] = 8'b01010101;
		data[164] = 8'b00111100;
		data[165] = 8'b00000010;
		data[166] = 8'b01011110;
		data[167] = 8'b11000110;
		data[168] = 8'b00110100;
		data[169] = 8'b01000010;
		data[170] = 8'b10010000;
		data[171] = 8'b10111101;
		data[172] = 8'b00000000;
		data[173] = 8'b00100010;
		data[174] = 8'b11111000;
		data[175] = 8'b00100101;
		// 1735311820 XOR 231278533 = 1789380105
		//H 676ec1cc XOR 0dc907c5 = 6aa7c609
		data[176] = 8'b00111100;
		data[177] = 8'b00000001;
		data[178] = 8'b01100111;
		data[179] = 8'b01101110;
		data[180] = 8'b00110100;
		data[181] = 8'b00100001;
		data[182] = 8'b11000001;
		data[183] = 8'b11001100;
		data[184] = 8'b00111100;
		data[185] = 8'b00000010;
		data[186] = 8'b00001101;
		data[187] = 8'b11001001;
		data[188] = 8'b00110100;
		data[189] = 8'b01000010;
		data[190] = 8'b00000111;
		data[191] = 8'b11000101;
		data[192] = 8'b00000000;
		data[193] = 8'b00100010;
		data[194] = 8'b11111000;
		data[195] = 8'b00100110;
		// 431714708 XORI 38687 = 431744651
		//H 19bb7194 XORI 0000971f = 19bbe68b
		data[196] = 8'b00111100;
		data[197] = 8'b00000001;
		data[198] = 8'b00011001;
		data[199] = 8'b10111011;
		data[200] = 8'b00110100;
		data[201] = 8'b00100001;
		data[202] = 8'b01110001;
		data[203] = 8'b10010100;
		data[204] = 8'b00111000;
		data[205] = 8'b00111111;
		data[206] = 8'b10010111;
		data[207] = 8'b00011111;
		// 1438218084 SLLV 3431212682 = 3359795360
		//H 55b97764 SLLV cc84268a = c84268a0
		data[208] = 8'b00111100;
		data[209] = 8'b00000001;
		data[210] = 8'b01010101;
		data[211] = 8'b10111001;
		data[212] = 8'b00110100;
		data[213] = 8'b00100001;
		data[214] = 8'b01110111;
		data[215] = 8'b01100100;
		data[216] = 8'b00111100;
		data[217] = 8'b00000010;
		data[218] = 8'b11001100;
		data[219] = 8'b10000100;
		data[220] = 8'b00110100;
		data[221] = 8'b01000010;
		data[222] = 8'b00100110;
		data[223] = 8'b10001010;
		data[224] = 8'b00000000;
		data[225] = 8'b00100010;
		data[226] = 8'b11111000;
		data[227] = 8'b00000100;
		// 3538836615 SLL 28 = 1879048192
		//H d2ee5c87 SLL 0000001c = 70000000
		data[228] = 8'b00111100;
		data[229] = 8'b00000001;
		data[230] = 8'b11010010;
		data[231] = 8'b11101110;
		data[232] = 8'b00110100;
		data[233] = 8'b00100001;
		data[234] = 8'b01011100;
		data[235] = 8'b10000111;
		data[236] = 8'b00000000;
		data[237] = 8'b00000001;
		data[238] = 8'b11111111;
		data[239] = 8'b00000000;
		// 2645139758 SRAV 811140775 = 49508
		//H 9da9a12e SRAV 305906a7 = 0000c164
		data[240] = 8'b00111100;
		data[241] = 8'b00000001;
		data[242] = 8'b10011101;
		data[243] = 8'b10101001;
		data[244] = 8'b00110100;
		data[245] = 8'b00100001;
		data[246] = 8'b10100001;
		data[247] = 8'b00101110;
		data[248] = 8'b00111100;
		data[249] = 8'b00000010;
		data[250] = 8'b00110000;
		data[251] = 8'b01011001;
		data[252] = 8'b00110100;
		data[253] = 8'b01000010;
		data[254] = 8'b00000110;
		data[255] = 8'b10100111;
		data[256] = 8'b00000000;
		data[257] = 8'b00100010;
		data[258] = 8'b11111000;
		data[259] = 8'b00000111;
		// 3986905438 SRA 4 = 1152921504587593109
		//H eda3595e SRA 00000004 = 0xfffffff_feda3595
		data[260] = 8'b00111100;
		data[261] = 8'b00000001;
		data[262] = 8'b11101101;
		data[263] = 8'b10100011;
		data[264] = 8'b00110100;
		data[265] = 8'b00100001;
		data[266] = 8'b01011001;
		data[267] = 8'b01011110;
		data[268] = 8'b00000000;
		data[269] = 8'b00000001;
		data[270] = 8'b11111001;
		data[271] = 8'b00000011;
		// 2538966711 SRLV 155967169 = 18
		//H 97558eb7 SRLV 094bdec1 = 00000012
		data[272] = 8'b00111100;
		data[273] = 8'b00000001;
		data[274] = 8'b10010111;
		data[275] = 8'b01010101;
		data[276] = 8'b00110100;
		data[277] = 8'b00100001;
		data[278] = 8'b10001110;
		data[279] = 8'b10110111;
		data[280] = 8'b00111100;
		data[281] = 8'b00000010;
		data[282] = 8'b00001001;
		data[283] = 8'b01001011;
		data[284] = 8'b00110100;
		data[285] = 8'b01000010;
		data[286] = 8'b11011110;
		data[287] = 8'b11000001;
		data[288] = 8'b00000000;
		data[289] = 8'b00100010;
		data[290] = 8'b11111000;
		data[291] = 8'b00000110;
		// 2052318909 SRL 16 = 31315
		//H 7a53e6bd SRL 00000010 = 00007a53
		data[292] = 8'b00111100;
		data[293] = 8'b00000001;
		data[294] = 8'b01111010;
		data[295] = 8'b01010011;
		data[296] = 8'b00110100;
		data[297] = 8'b00100001;
		data[298] = 8'b11100110;
		data[299] = 8'b10111101;
		data[300] = 8'b00000000;
		data[301] = 8'b00000001;
		data[302] = 8'b11111100;
		data[303] = 8'b00000010;
	end
endmodule

module Memory(clk, rw_mem, mem_ref,
			  mem_addr, din, dout);
	input clk;
	input rw_mem;
	input [31:0] mem_addr;
	input [7:0] din;

	output reg mem_ref;
	output reg [7:0] dout;

    reg [7:0] data[1023:0];
	
	always @(negedge clk)
	begin
		if (rw_mem == `READ_VALID)
		begin
			dout = data[mem_addr];
			mem_ref = `FULL;
		end
		else if (rw_mem == `WRITE_VALID)
		begin
			data[mem_addr] = din;
			mem_ref = `FULL;
		end
		else
		begin
			mem_ref = `EMPTY;
		end
	end

endmodule